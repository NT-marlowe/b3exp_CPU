`include "define.vh"

module alu(
    input wire [5:0] alucode,
    input wire [31:0] op1,
    input wire [31:0] op2,
    output reg [31:0] alu_result,
    output reg br_taken // 分岐の有無
);

    // always @(alucode or op1 or op2) begin
    always @(*) begin
        case (alucode) 
            `ALU_LUI : begin
                alu_result <= op2;
                br_taken <= `DISABLE;
            end

            `ALU_JAL : begin
                alu_result <= op2 + 3'd4;
                br_taken <= `ENABLE;
            end

            `ALU_JALR : begin
                alu_result <= op2 + 3'd4;
                br_taken <= `ENABLE;
            end

            `ALU_BEQ : begin
                alu_result <= 1'b0;
                br_taken <= (op1 == op2)? `ENABLE : `DISABLE;
            end

            `ALU_BNE : begin
                alu_result <= 1'b0;
                br_taken <= (op1 != op2)? `ENABLE : `DISABLE;
            end

            `ALU_BLT : begin
                alu_result <= 1'b0;
                br_taken <= ($signed(op1) < $signed(op2))? `ENABLE : `DISABLE;
            end

            `ALU_BGE : begin
                alu_result <= 1'b0;
                br_taken <= ($signed(op1) >= $signed(op2))? `ENABLE : `DISABLE;
            end

            `ALU_BLTU : begin
                alu_result <= 1'b0;
                br_taken <= (op1 < op2)? `ENABLE : `DISABLE;
            end

            `ALU_BGEU : begin
                alu_result <= 1'b0;
                br_taken <= (op1 >= op2)? `ENABLE : `DISABLE;
            end

            `ALU_LB, `ALU_LH, `ALU_LW, `ALU_LBU, `ALU_LHU : begin
                alu_result <= op1 + op2;
                br_taken <= `DISABLE;
            end

            // `ALU_LW : begin
            //     alu_result <= op1 + op2;
            //     br_taken <= `DISABLE;
            // end

            // `ALU_LBU : begin
            //     alu_result <= op1 + op2;
            //     br_taken <= `DISABLE
            // end

            // `ALU_LHU : begin
            //     alu_result <= op1 + op2;
            //     br_taken <= `DISABLE
            // end

            `ALU_SB, `ALU_SH, `ALU_SW : begin
                alu_result <= op1 + op2;
                br_taken <= `DISABLE;
            end

            // `ALU_SH : begin
            //     alu_result <= op1 + op2;
            //     br_taken <= `DISABLE;
            // end

            // `ALU_SW : begin
            //     alu_result <= op1 + op2;
            //     br_taken <= `DISABLE;
            // end

            `ALU_ADD : begin
                alu_result <= op1 + op2;
                br_taken <= `DISABLE;
            end

            `ALU_SUB : begin
                alu_result <= op1 - op2;
                br_taken <= `DISABLE;
            end

            `ALU_SLT :begin
                alu_result <= ($signed(op1) < $signed(op2))? 1'b1 : 1'b0;
                br_taken <= `DISABLE;
            end

            `ALU_SLTU : begin 
                alu_result <= (op1 < op2)? 1'b1 : 1'b0;
                br_taken <= `DISABLE;
            end

            `ALU_XOR : begin
                alu_result <= op1 ^ op2;
                br_taken <= `DISABLE;
            end

            `ALU_OR : begin
                alu_result <= op1 | op2;
                br_taken <= `DISABLE;
            end
            
            `ALU_AND : begin
                alu_result <= op1 & op2;
                br_taken <= `DISABLE;
            end

            `ALU_SLL : begin 
                alu_result <= op1 << op2[4:0];
                br_taken <= `DISABLE;
            end

            `ALU_SRL : begin
                alu_result <= op1 >> op2[4:0];
                br_taken <= `DISABLE;
            end

            `ALU_SRA : begin
                alu_result <= ($signed(op1) >>> op2[4:0]);
                br_taken <= `DISABLE;
            end

            `ALU_NOP : begin
                alu_result <= 1'b0;
                br_taken <= `DISABLE;
            end

            default : begin
                alu_result <= 1'b0;
                br_taken <= `DISABLE;
            end
        endcase
    end

endmodule